module Mcu_tb; 
    reg clk, reset,
    


endmodule