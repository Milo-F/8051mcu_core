/*----------------------------------------
 *    File Name: IntArbiter.v
 *    function: Interupt arbiter to orgnize the priority of interupt
 *    author: Milo
 *    Data: 2022-02-24
 *    Version: 1.0
----------------------------------------*/

module IntArbiter(
    input int0,
    input int1,
    input t0,
    input t1,
    input uart,
    // output
    output int_early
);

endmodule