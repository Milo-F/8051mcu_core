module Timer(
    input clk,
    input rst_n,
    input[7:0] tcon_in, tmod_in, tl0_in, tl1_in, th0_in, th1_in,
    output[7:0] tcon_out, tmod_out, tl0_out, tl1_out, th0_out, th1_out
);

endmodule