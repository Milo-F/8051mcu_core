module UartCtl (
    input                   clk,
    input                   rst_n,
    
);

endmodule