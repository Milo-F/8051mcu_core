module FullAdder (
    a, b, c_in, sum, c_out
);
    input a, b, c_in;
    output sum, c_out;
    
endmodule