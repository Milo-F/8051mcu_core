/*----------------------------------------
 *    File Name: rtl/UartIf.v
 *    function: Uart interface, transmite the data from fifo, and receive the data to fifo.
 *    author: Milo
 *    Data: 2022-03-10
 *    Version: 1.0
 ----------------------------------------*/

module UartIf (
    input                                                   clk_uart,
    input                                                   rst_n,
    input                   [7:0]                           txd_from_fifo,
    input                                                   fifo_empty,    // if fifo is empty, stop transimiting
    output                                                  r_en,
    output                                                  txd,
    input                                                   rxd_int_in,    // 接收中断标志位
    input                                                   rxd,
    output                  [7:0]                           r_data,
    output                                                  rxd_int
);
    /*
     *   串口发送
     */
    wire                    clk_tx; // 发送时钟，波特率9600
    reg                     clk_rd; // 读fifo时钟，发送时钟的12分频，包括1起始位+8数据位+1校验位+2空闲位
    reg         [3:0]       tx_bit_cnt, tx_bit_cnt_nxt; // 发送数据计数，记录已经发了几个bit
    reg                     txd_out, txd_out_nxt;
    reg                     tx_status, tx_status_nxt;
    reg         [11:0]      tx_tmp, tx_tmp_nxt;
    wire                    odd_bit;
    wire        [3:0]       tx_bit_cnt_minus_1;
    
    assign tx_bit_cnt_minus_1 = tx_bit_cnt - 1;
    assign odd_bit            = ^txd_from_fifo;
    assign txd                = txd_out;
    // wire clk_tx;
    ClkDiv #(
        .DIV_NUM(16)
    ) ClkDiv_tx (
        .clk_in(clk_uart),
        .rst_n(rst_n),
        .clk_out(clk_tx)
    );
    
    always @* begin
        tx_bit_cnt_nxt = 4'b1011;
        clk_rd         = 0;
        tx_status_nxt  = 0;
        if (!fif o_empty) begin
            tx_status_nxt = 1;
            if (tx_bit_cnt == 0) begin
                tx_bit_cnt_nxt = 4'b1011;
                clk_rd         = 1;
            end
            else begin
                tx_bit_cnt_nxt = tx_bit_cnt_minus_1;
            end
        end
    end
    
    assign r_en = clk_rd; // 按照读时钟去读数据
    
    always @* begin
        txd_out_nxt   = 1;
        tx_tmp_nxt    = tx_tmp;
        tx_status_nxt = tx_status;
        
        if (tx_status) begin // 发送数据
            txd_out_nxt = tx_tmp[0];
            tx_tmp_nxt  = {1, tx_tmp[11:1]};
        end
    end
    
    always @(posedge clk_tx) begin
        if (!rst_n) begin
            tx_status  <= 0;
            txd_out    <= 1;
            tx_tmp     <= 12'hfff;
            tx_bit_cnt <= 4'b1011;
        end
        else begin
            tx_status  <= tx_status_nxt;
            txd_out    <= txd_out_nxt;
            tx_tmp     <= r_en ? {2'b11, odd_bit, txd_from_fifo, 1'b0} : tx_tmp_nxt;
            tx_bit_cnt <= tx_bit_cnt_nxt;
        end
    end
    /*
     *   串口接收：串口接收16倍波特率采样，波特率9600
     */
    // 计数器等寄存器声明
    reg                     int_hold, int_hold_nxt; // 中断保持
    reg         [7:0]       r_data_out, r_data_out_nxt;
    reg                     rxd_int_out, rxd_int_out_nxt;
    reg         [8:0]       rx_tmp, rx_tmp_nxt;
    reg                     rx_status, rx_status_nxt; // 0 : wait  1 : busy
    reg         [2:0]       start_cnt, start_cnt_nxt;
    reg         [3:0]       sample_cnt, sample_cnt_nxt;
    reg         [3:0]       bit_cnt, bit_cnt_nxt;
    wire        [2:0]       start_cnt_minus_1;
    wire        [3:0]       sample_cnt_minus_1;
    wire        [3:0]       bit_cnt_minus_1;
    // counter
    assign start_cnt_minus_1  = start_cnt - 1;
    assign sample_cnt_minus_1 = sample_cnt - 1;
    assign bit_cnt_minus_1    = bit_cnt - 1;
    // receive out
    assign rxd_int = rxd_int_out;
    assign r_data  = r_data_out;
    
    // 串口接收组合逻辑
    always @* begin
        int_hold_nxt    = rxd_int_in ? 1'b0 : int_hold; // 等到中断标志为1再取消保持
        r_data_out_nxt  = r_data_out;
        rxd_int_out_nxt = (int_hold) ? rxd_int_out : rxd_int_in; // 接收中断需要持续大于等于两个周期
        start_cnt_nxt   = start_cnt;
        sample_cnt_nxt  = sample_cnt;
        rx_status_nxt   = rx_status;
        bit_cnt_nxt     = bit_cnt;
        rx_tmp_nxt      = rx_tmp;
        if (!rx_status) begin // when bus is empty : detecting 0
            if (!rxd) begin
                if (start_cnt == 3'b0) begin
                    rx_status_nxt  = 1;
                    bit_cnt_nxt    = 4'b1010;
                    sample_cnt_nxt = 3'b111;
                end
                start_cnt_nxt = start_cnt_minus_1;
            end
            else begin
                start_cnt_nxt = 4'b1111;
            end
        end
        else begin
            sample_cnt_nxt = sample_cnt_minus_1;
            if (sample_cnt == 4'b0) begin // sample
                rx_tmp_nxt  = {rxd, rx_tmp[8:1]};
                bit_cnt_nxt = bit_cnt_minus_1;
            end
            
            if (bit_cnt == 4'b0) begin
                rx_status_nxt   = 0;
                rxd_int_out_nxt = 1'b1;
                rx_tmp_nxt      = 9'b0;
                int_hold_nxt    = ~rxd_int;
                // 奇校验
                r_data_out_nxt = rx_tmp[8] == (^rx_tmp[7:0]) ? rx_tmp[7:0] : 8'b0;
            end
        end
    end
    // 次态传递
    always @(posedge clk_uart) begin
        if (!rst_n) begin
            r_data_out  <= 0;
            rxd_int_out <= 0;
            start_cnt   <= 3'b111;
            sample_cnt  <= 4'b1111;
            bit_cnt     <= 4'b1010;
            rx_status   <= 0;
            rx_tmp      <= 0;
            int_hold    <= 0;
        end
        else begin
            int_hold    <= int_hold_nxt;
            r_data_out  <= r_data_out_nxt;
            rxd_int_out <= rxd_int_out_nxt;
            start_cnt   <= start_cnt_nxt;
            sample_cnt  <= sample_cnt_nxt;
            bit_cnt     <= bit_cnt_nxt;
            rx_status   <= !rxd_int_in & rx_status_nxt; // must solve the interupt to continue receiv data
            rx_tmp      <= rx_tmp_nxt;
        end
    end
endmodule
