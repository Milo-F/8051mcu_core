module top_tb_mcu();
    
endmodule